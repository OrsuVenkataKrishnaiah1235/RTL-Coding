module Ripple_Carry_Adder
