module top_module ( input a, input b, output out );
    mod_a hi(a,b,out);
endmodule